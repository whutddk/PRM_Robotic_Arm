module prm_oblgc_chk630
(
input A,
input B,
input C,
input D,
input E,
input F,
input G,
input H,
input I,
input J,
input K,
input L,
input M,
input N,
input O,
output edge_mask
);
assign edge_mask = (!O&N&M&!J&I&H&G&F&E&!D)|(!O&M&!L&!K&!J&I&H&F&!E&D&B&A)|(!O&N&L&J&!I&!H&!G&D&!C&!B&!A)|(!O&N&L&K&J&!I&!H&!G&!F&D&!C&!B)|(N&!M&K&!J&I&H&G&!E&D&A)|(!O&N&M&!J&I&H&G&!E&C&B&A)|(!N&M&K&!J&I&H&G&F&E&!D&!B&!A)|(!L&K&!J&I&H&G&F&!E&D&B&A)|(!M&L&!J&I&H&G&!E&D&!C&B&A)|(O&!N&!L&!K&!J&I&H&F&!E&D&!A)|(O&!M&!L&!K&!J&I&H&G&!D&C&!B&!A)|(!M&!L&K&J&!I&!H&!F&!E&D&C&!B&!A)|(!L&!K&J&!I&!H&!G&!E&D&B&!A)|(O&!N&!L&!J&I&H&G&F&E&!D)|(!M&L&K&!J&I&H&G&F&E&!D&!C&!A)|(!M&L&J&!I&!H&!G&!F&E&!D&!C)|(!M&L&K&!J&I&H&G&E&!D&!C&!B&!A)|(O&!N&!K&J&!I&!H&!G&!F&D&!C&!B&!A)|(N&!M&L&K&J&!I&!H&!F&!E&D&!A)|(N&!M&!J&I&H&G&F&E&!D&!B&!A)|(O&!N&!M&J&!I&!H&!G&!F&D&!C&!B)|(!M&L&K&J&!I&!H&!G&E&!D&!C)|(!M&L&K&J&!I&!H&!G&!E&D&B)|(O&!K&!J&I&H&G&F&!E&C&B)|(!O&!N&!M&L&J&!I&!H&!F&E&!D&!C&!B&A)|(O&!N&!L&!K&J&!I&!H&!F&!E&D&!A)|(O&!N&M&!L&!K&J&!I&!H&!F&!D&C&B&!A)|(O&!K&J&!I&!H&!G&!E&!D&C&B&A)|(O&!N&!L&K&J&!I&!H&!F&E&!D&C&!B)|(O&!L&K&J&!I&!H&!G&!F&!E&B&A)|(O&!K&J&!I&!H&!G&!F&!E&C&B)|(O&!M&!J&I&H&G&!E&C&B)|(O&!M&L&J&!I&!H&!F&!E&D)|(O&!M&!L&J&!I&!H&!G&!F&!E)|(N&!M&!L&!K&!J&I&H&G&F&E&!D&!A)|(!O&N&K&J&!I&!H&!F&!E&D&!C&A)|(!M&L&!J&I&H&G&!E&D&C&!B)|(O&!N&!K&!J&I&H&G&F&E&!D)|(!N&M&K&!J&I&H&G&E&!D&!C)|(O&N&!L&!K&!J&I&H&G&F&!D&!C&B&!A)|(!N&M&L&K&!J&I&H&G&E&!D&!B&!A)|(!N&M&L&K&J&!I&!H&!G&E&!D)|(O&L&!K&!J&I&H&G&F&!E&C&A)|(O&!M&!K&!J&I&H&G&!D&!C&B&!A)|(!O&!N&M&L&J&!I&!H&!F&E&!D&C&!B&A)|(O&!N&!M&J&!I&!H&!G&D&!C&!B&!A)|(O&!N&M&!K&J&!I&!H&!F&E&!D&C&!B)|(N&M&!L&!K&J&!I&!H&!F&!E&D&!C)|(O&!N&!M&!J&I&H&G&!D&C&B&!A)|(O&!N&!M&!J&I&H&G&F&E&!D)|(O&N&!L&!J&I&H&G&F&!E&B&A)|(O&!N&L&!K&!J&I&H&G&!E&B)|(O&!M&!K&J&!I&!H&!G&!F&!E)|(!O&N&M&!J&I&H&G&F&D&!C&!B&!A)|(O&!M&!K&J&!I&!H&!G&!E&B)|(!O&N&L&K&!J&I&H&F&!E&D&!A)|(O&!N&M&L&!J&I&H&G&!E&C)|(O&!N&!M&L&J&!I&!H&!F&!D&C&B&!A)|(!O&N&L&!J&I&H&F&!E&D&!C)|(O&N&!M&J&!I&!H&!G&!F&!E&B)|(!N&!M&L&K&!J&I&H&F&!E&D&C)|(O&!N&J&!I&!H&!G&!E&C&B)|(!L&K&!J&I&H&G&F&!E&D&C)|(O&!N&M&L&J&!I&!H&!G&!F&!D)|(!M&L&K&!J&I&H&G&F&E&!D&!C&!B)|(M&!L&!K&J&!I&!H&!G&E&!D&!C&!A)|(!M&L&!J&I&H&G&!E&D&C&!A)|(!N&!M&L&!J&I&H&F&!E&D&!C&B&A)|(O&L&!K&J&!I&!H&!G&!F&!E&C&A)|(O&!N&!M&!J&I&H&G&F&D&!C&!B&!A)|(O&!K&!J&I&H&G&F&!E&D)|(!N&M&!J&I&H&G&F&E&!D&!C)|(!N&M&K&J&!I&!H&!G&E&!D&!A)|(O&!M&!L&!J&I&H&G&!E&A)|(!N&M&!J&I&H&G&E&!D&!C&!B)|(!M&J&!I&!H&!G&!E&D&!C&B&A)|(O&!N&!L&!J&I&H&F&!E&D&!B)|(O&!L&J&!I&!H&!G&!E&D)|(!N&M&!K&J&!I&!H&!F&E&!D&C&!B&!A)|(O&!N&!L&J&!I&!H&!G&D&!C&!B&!A)|(M&!L&!J&I&H&G&F&E&!D&!C&!B)|(N&M&!L&J&!I&!H&!G&!E&C&B&A)|(N&M&!L&!K&J&!I&!H&!F&!E&D&!B)|(O&N&!L&!K&J&!I&!H&!G&!F&!D&!C&B)|(O&!N&!L&!J&I&H&G&E&!D&!A)|(!N&M&!L&K&J&!I&!H&!F&E&!D&C&!B)|(O&!N&K&J&!I&!H&!F&E&!D&C&!B&!A)|(O&N&!M&J&!I&!H&!G&!F&!E&A)|(O&!N&M&K&J&!I&!H&!G&!D&C)|(O&!N&!M&L&J&!I&!H&!F&E&!D&C&!B)|(N&!L&K&J&!I&!H&!G&!E&D&A)|(N&!M&!J&I&H&G&!E&D&C)|(!M&L&!J&I&H&G&F&E&!D&!C&!B&!A)|(!M&L&K&!J&I&H&G&!E&D&B)|(O&N&!M&!J&I&H&G&F&!E&A)|(!M&L&K&J&!I&!H&!G&E&!D&!B&!A)|(O&!M&!L&!J&I&H&G&F&!D&!B)|(!N&M&J&!I&!H&!G&E&!D&!C)|(!O&N&M&K&J&!I&!H&!G&!D)|(!N&M&L&!J&I&H&G&F&E&!D&!B)|(N&!L&J&!I&!H&!G&E&!D&!C&!B)|(O&!N&!K&!J&I&H&G&E&!D&!B)|(!N&M&L&J&!I&!H&!G&E&!D&!A)|(N&!M&!J&I&H&G&E&!D&!C&!B)|(O&!M&!L&!J&I&H&G&!D&!C&B)|(O&!N&!L&K&!J&I&H&G&!D&C&!B)|(O&!N&!L&K&!J&I&H&G&!E&A)|(O&!M&!L&J&!I&!H&!G&!E&A)|(O&!N&M&K&!J&I&H&G&!E&B)|(O&!N&L&!K&J&!I&!H&!G&!D&C)|(O&!N&M&K&J&!I&!H&!G&!D&A)|(!O&!M&L&!J&I&H&F&!E&D&C&!B)|(O&!L&!J&I&H&G&!E&D&!B&!A)|(!N&M&!J&I&H&G&!E&D&C)|(O&!M&!K&!J&I&H&G&F&!D&!B)|(!N&M&J&!I&!H&!G&!E&D&B)|(N&!M&L&J&!I&!H&!F&!E&D&!C)|(!N&M&L&!J&I&H&G&E&!D&!C)|(O&!L&!J&I&H&G&!E&D&!C)|(!M&L&J&!I&!H&!G&E&!D&!C&!B)|(N&!M&L&J&!I&!H&!G&!E&D)|(O&N&!M&!J&I&H&G&F&!D&!C&B)|(O&!N&M&L&!J&I&H&G&F&!D&!A)|(O&!M&!L&J&!I&!H&!G&!D&C&!B)|(O&N&!M&J&!I&!H&!G&!D&!C&B&A)|(O&!N&L&!K&J&!I&!H&!G&!D&A)|(O&!N&M&L&!J&I&H&G&!E&A)|(O&!N&!L&K&J&!I&!H&!G&!D&B)|(!K&J&!I&!H&!G&!E&D&C&!B)|(L&!K&!J&I&H&G&F&!E&D&B)|(!O&N&M&!J&I&H&G&!E&D)|(!O&N&M&J&!I&!H&!G&D&!C&!B)|(O&!N&M&L&J&!I&!H&!G&!D&B)|(N&!M&!J&I&H&G&!E&D&B)|(!O&N&M&L&J&!I&!H&!G&!E)|(!N&M&!J&I&H&G&!E&D&B)|(!L&K&J&!I&!H&!G&E&!D&!C&!B)|(!N&J&!I&!H&!G&!F&!E&D&B)|(N&!M&L&J&!I&!H&!F&!E&D&!B)|(O&!K&J&!I&!H&!G&!E&D&!C)|(!M&L&J&!I&!H&!G&E&!D&!C&!A)|(!N&M&J&!I&!H&!G&E&!D&!B)|(O&!M&!K&J&!I&!H&!G&!D&C&!B)|(O&!M&!L&J&!I&!H&!G&!D&B&!A)|(!K&J&!I&!H&!G&!E&D&C&!A)|(!L&K&J&!I&!H&!G&!E&D&C)|(!O&L&J&!I&!H&!G&!E&D&C)|(N&!L&J&!I&!H&!G&!E&D&B)|(N&!M&L&!J&I&H&G&!E&D)|(!O&N&L&!J&I&H&G&F&E&!D)|(!O&N&K&!J&I&H&G&F&E&!D)|(!O&N&!J&I&H&G&E&!D&!B)|(!O&N&M&L&!J&I&H&G&!D)|(!O&N&M&K&!J&I&H&G&!D)|(!O&N&M&!J&I&H&G&E&!D&!A)|(!O&N&!J&I&H&G&E&!D&!C)|(!O&N&L&!J&I&H&G&E&!D&!A)|(!O&!N&M&!J&I&H&F&E&!D&!C&!B)|(!O&!N&M&L&!K&!J&I&H&F&E&!D&!C&!A)|(!O&!N&M&!L&K&!J&I&H&F&E&!D&!C&!A)|(!O&!N&L&K&!J&I&H&F&E&!D&!C&!B&!A)|(O&!N&!M&!J&I&H&G&E&!D&!B)|(O&!N&!M&!L&!J&I&H&G&!D)|(O&!N&!M&!K&!J&I&H&G&!D)|(O&!N&!J&I&H&G&E&!D&!C)|(!O&N&M&J&!I&!H&!F&D&!C&!B&!A)|(!O&N&L&J&!I&!H&!F&D&!C&!B&!A)|(!O&N&K&J&!I&!H&!G&E&!C&!B&!A)|(!O&N&!M&J&!I&!H&!F&E&!D&C&B&A)|(!N&M&!L&J&!I&!H&!F&E&!D&!C&B&A)|(!O&!N&M&L&J&!I&!H&!F&E&!D&C&B&!A)|(!O&!N&!M&L&!K&J&!I&!H&!F&E&!D&!C&!B)|(!O&N&J&!I&!H&!G&E&!D)|(!O&N&!M&!L&J&!I&!H&!F&E&!D&C&B)|(!O&!N&M&!L&!K&J&!I&!H&!F&E&!D&!C&B)|(!O&!N&!M&L&K&J&!I&!H&!F&E&!D&!C&B)|(!O&M&!L&!J&I&H&F&!E&D&C)|(!O&M&!K&!J&I&H&F&!E&D&C&B&A)|(!O&N&M&!J&I&H&F&!E&D)|(!N&!M&L&!J&I&H&F&!E&D&C&!A)|(!O&N&K&!J&I&H&F&!E&D&!C&A)|(!O&N&K&!J&I&H&F&!E&D&C&!B&!A)|(!O&N&!J&I&H&F&!E&D&!C&B&!A)|(O&!N&!M&!L&J&!I&!H&!F&D&!C&!B&!A)|(O&!N&!M&!K&J&!I&!H&!G&!C&!B)|(O&!N&!M&!L&J&!I&!H&!G&!C&!B)|(!O&N&M&!J&I&H&F&!E&C&B&A)|(!O&N&M&L&!J&I&H&F&!E)|(!O&N&M&K&!J&I&H&F&!E)|(O&!N&M&L&J&!I&!H&!F&E&!D&!C&B)|(O&!N&!J&I&H&G&!E&D)|(O&!N&M&L&K&J&!I&!H&!F&E&!D&!C)|(O&!N&J&!I&!H&!G&E&!D)|(O&N&!M&!L&!K&J&!I&!H&!F&E&!D&!C)|(O&!N&M&K&J&!I&!H&!F&E&!D&!C&B)|(O&N&!M&!K&J&!I&!H&!F&E&!D&!C&!B)|(O&N&!M&!L&J&!I&!H&!F&E&!D&!C&!B)|(O&N&!M&!L&J&!I&!H&!F&E&!D&!C&!A)|(O&N&!M&J&!I&!H&!F&E&!D&!C&!B&!A)|(O&!N&!K&!J&I&H&F&!E&D&!C)|(O&!N&!L&!J&I&H&F&!E&D&!C)|(O&!N&!K&!J&I&H&F&!E&D&!B&!A)|(O&!N&!J&I&H&F&!E&D&!C&!B)|(O&!N&!J&I&H&F&!E&D&!C&!A)|(O&!N&!J&I&H&F&!E&!D&C&B)|(O&!L&!K&!J&I&H&G&!E&C&B)|(O&N&!L&!J&I&H&G&F&!E&C)|(O&N&!M&!J&I&H&G&!E&C)|(O&N&!L&!K&!J&I&H&G&!E&C&A)|(O&!N&!M&!K&!J&I&H&F&!E)|(O&!N&!M&!L&!J&I&H&F&!E)|(O&N&!M&!J&I&H&G&!E&B&A)|(!N&!M&L&!K&J&!I&!H&!F&!E&D&C&B&A)|(!N&!M&!L&K&J&!I&!H&!F&!E&D&C)|(!O&N&M&J&!I&!H&!F&!E&D)|(!N&!M&!L&J&!I&!H&!F&!E&D&!C&B&A)|(!O&N&J&!I&!H&!F&!E&D&!C&B&!A)|(!O&N&M&J&!I&!H&!F&!E&C&B&A)|(!O&N&M&L&J&!I&!H&!F&!E)|(!O&N&M&K&J&!I&!H&!F&!E)|(O&!N&!L&J&!I&!H&!F&!E&D&!B)|(O&!M&J&!I&!H&!F&!E&D&C&B&A)|(O&!N&!K&J&!I&!H&!F&!E&D&!C)|(O&!N&!L&J&!I&!H&!F&!E&D&!C)|(O&!N&!K&J&!I&!H&!F&!E&D&!B&!A)|(O&!M&K&J&!I&!H&!F&!E&D&!B)|(O&!N&J&!I&!H&!F&!E&D&!C&!B)|(O&!M&L&J&!I&!H&!F&!E&C&B)|(O&!M&K&J&!I&!H&!F&!E&C&B)|(O&!N&J&!I&!H&!F&!E&D&!C&!A)|(O&!N&J&!I&!H&!G&!E&D)|(O&!N&J&!I&!H&!F&!E&!D&C&B)|(O&!N&!M&!K&J&!I&!H&!F&!E)|(O&N&!M&L&J&!I&!H&!F&!E&C&A)|(O&!N&!M&!L&J&!I&!H&!F&!E)|(O&N&!L&!K&J&!I&!H&!G&!E&C&A)|(O&N&!M&J&!I&!H&!G&!E&C)|(O&!L&!K&J&!I&!H&!G&!E&C&B)|(O&N&!L&J&!I&!H&!G&!F&!E&C);
endmodule