module prm_lgcchk_top
(
input A,
input B,
input C,
input D,
input E,
input F,
input G,
input H,
input I,
input J,
input K,
input L,
input M,
input N,
input O,
output [1023:0] edge_mask
);
prm_oblgc_chk0 i_prm_oblgc_chk0(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[0])
);
prm_oblgc_chk1 i_prm_oblgc_chk1(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1])
);
prm_oblgc_chk2 i_prm_oblgc_chk2(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[2])
);
prm_oblgc_chk3 i_prm_oblgc_chk3(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[3])
);
prm_oblgc_chk4 i_prm_oblgc_chk4(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[4])
);
prm_oblgc_chk5 i_prm_oblgc_chk5(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[5])
);
prm_oblgc_chk6 i_prm_oblgc_chk6(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[6])
);
prm_oblgc_chk7 i_prm_oblgc_chk7(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[7])
);
prm_oblgc_chk8 i_prm_oblgc_chk8(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[8])
);
prm_oblgc_chk9 i_prm_oblgc_chk9(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[9])
);
prm_oblgc_chk10 i_prm_oblgc_chk10(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[10])
);
prm_oblgc_chk11 i_prm_oblgc_chk11(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[11])
);
prm_oblgc_chk12 i_prm_oblgc_chk12(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[12])
);
prm_oblgc_chk13 i_prm_oblgc_chk13(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[13])
);
prm_oblgc_chk14 i_prm_oblgc_chk14(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[14])
);
prm_oblgc_chk15 i_prm_oblgc_chk15(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[15])
);
prm_oblgc_chk16 i_prm_oblgc_chk16(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[16])
);
prm_oblgc_chk17 i_prm_oblgc_chk17(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[17])
);
prm_oblgc_chk18 i_prm_oblgc_chk18(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[18])
);
prm_oblgc_chk19 i_prm_oblgc_chk19(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[19])
);
prm_oblgc_chk20 i_prm_oblgc_chk20(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[20])
);
prm_oblgc_chk21 i_prm_oblgc_chk21(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[21])
);
prm_oblgc_chk22 i_prm_oblgc_chk22(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[22])
);
prm_oblgc_chk23 i_prm_oblgc_chk23(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[23])
);
prm_oblgc_chk24 i_prm_oblgc_chk24(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[24])
);
prm_oblgc_chk25 i_prm_oblgc_chk25(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[25])
);
prm_oblgc_chk26 i_prm_oblgc_chk26(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[26])
);
prm_oblgc_chk27 i_prm_oblgc_chk27(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[27])
);
prm_oblgc_chk28 i_prm_oblgc_chk28(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[28])
);
prm_oblgc_chk29 i_prm_oblgc_chk29(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[29])
);
prm_oblgc_chk30 i_prm_oblgc_chk30(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[30])
);
prm_oblgc_chk31 i_prm_oblgc_chk31(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[31])
);
prm_oblgc_chk32 i_prm_oblgc_chk32(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[32])
);
prm_oblgc_chk33 i_prm_oblgc_chk33(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[33])
);
prm_oblgc_chk34 i_prm_oblgc_chk34(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[34])
);
prm_oblgc_chk35 i_prm_oblgc_chk35(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[35])
);
prm_oblgc_chk36 i_prm_oblgc_chk36(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[36])
);
prm_oblgc_chk37 i_prm_oblgc_chk37(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[37])
);
prm_oblgc_chk38 i_prm_oblgc_chk38(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[38])
);
prm_oblgc_chk39 i_prm_oblgc_chk39(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[39])
);
prm_oblgc_chk40 i_prm_oblgc_chk40(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[40])
);
prm_oblgc_chk41 i_prm_oblgc_chk41(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[41])
);
prm_oblgc_chk42 i_prm_oblgc_chk42(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[42])
);
prm_oblgc_chk43 i_prm_oblgc_chk43(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[43])
);
prm_oblgc_chk44 i_prm_oblgc_chk44(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[44])
);
prm_oblgc_chk45 i_prm_oblgc_chk45(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[45])
);
prm_oblgc_chk46 i_prm_oblgc_chk46(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[46])
);
prm_oblgc_chk47 i_prm_oblgc_chk47(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[47])
);
prm_oblgc_chk48 i_prm_oblgc_chk48(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[48])
);
prm_oblgc_chk49 i_prm_oblgc_chk49(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[49])
);
prm_oblgc_chk50 i_prm_oblgc_chk50(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[50])
);
prm_oblgc_chk51 i_prm_oblgc_chk51(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[51])
);
prm_oblgc_chk52 i_prm_oblgc_chk52(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[52])
);
prm_oblgc_chk53 i_prm_oblgc_chk53(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[53])
);
prm_oblgc_chk54 i_prm_oblgc_chk54(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[54])
);
prm_oblgc_chk55 i_prm_oblgc_chk55(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[55])
);
prm_oblgc_chk56 i_prm_oblgc_chk56(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[56])
);
prm_oblgc_chk57 i_prm_oblgc_chk57(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[57])
);
prm_oblgc_chk58 i_prm_oblgc_chk58(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[58])
);
prm_oblgc_chk59 i_prm_oblgc_chk59(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[59])
);
prm_oblgc_chk60 i_prm_oblgc_chk60(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[60])
);
prm_oblgc_chk61 i_prm_oblgc_chk61(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[61])
);
prm_oblgc_chk62 i_prm_oblgc_chk62(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[62])
);
prm_oblgc_chk63 i_prm_oblgc_chk63(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[63])
);
prm_oblgc_chk64 i_prm_oblgc_chk64(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[64])
);
prm_oblgc_chk65 i_prm_oblgc_chk65(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[65])
);
prm_oblgc_chk66 i_prm_oblgc_chk66(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[66])
);
prm_oblgc_chk67 i_prm_oblgc_chk67(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[67])
);
prm_oblgc_chk68 i_prm_oblgc_chk68(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[68])
);
prm_oblgc_chk69 i_prm_oblgc_chk69(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[69])
);
prm_oblgc_chk70 i_prm_oblgc_chk70(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[70])
);
prm_oblgc_chk71 i_prm_oblgc_chk71(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[71])
);
prm_oblgc_chk72 i_prm_oblgc_chk72(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[72])
);
prm_oblgc_chk73 i_prm_oblgc_chk73(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[73])
);
prm_oblgc_chk74 i_prm_oblgc_chk74(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[74])
);
prm_oblgc_chk75 i_prm_oblgc_chk75(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[75])
);
prm_oblgc_chk76 i_prm_oblgc_chk76(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[76])
);
prm_oblgc_chk77 i_prm_oblgc_chk77(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[77])
);
prm_oblgc_chk78 i_prm_oblgc_chk78(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[78])
);
prm_oblgc_chk79 i_prm_oblgc_chk79(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[79])
);
prm_oblgc_chk80 i_prm_oblgc_chk80(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[80])
);
prm_oblgc_chk81 i_prm_oblgc_chk81(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[81])
);
prm_oblgc_chk82 i_prm_oblgc_chk82(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[82])
);
prm_oblgc_chk83 i_prm_oblgc_chk83(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[83])
);
prm_oblgc_chk84 i_prm_oblgc_chk84(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[84])
);
prm_oblgc_chk85 i_prm_oblgc_chk85(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[85])
);
prm_oblgc_chk86 i_prm_oblgc_chk86(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[86])
);
prm_oblgc_chk87 i_prm_oblgc_chk87(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[87])
);
prm_oblgc_chk88 i_prm_oblgc_chk88(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[88])
);
prm_oblgc_chk89 i_prm_oblgc_chk89(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[89])
);
prm_oblgc_chk90 i_prm_oblgc_chk90(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[90])
);
prm_oblgc_chk91 i_prm_oblgc_chk91(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[91])
);
prm_oblgc_chk92 i_prm_oblgc_chk92(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[92])
);
prm_oblgc_chk93 i_prm_oblgc_chk93(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[93])
);
prm_oblgc_chk94 i_prm_oblgc_chk94(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[94])
);
prm_oblgc_chk95 i_prm_oblgc_chk95(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[95])
);
prm_oblgc_chk96 i_prm_oblgc_chk96(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[96])
);
prm_oblgc_chk97 i_prm_oblgc_chk97(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[97])
);
prm_oblgc_chk98 i_prm_oblgc_chk98(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[98])
);
prm_oblgc_chk99 i_prm_oblgc_chk99(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[99])
);
prm_oblgc_chk100 i_prm_oblgc_chk100(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[100])
);
prm_oblgc_chk101 i_prm_oblgc_chk101(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[101])
);
prm_oblgc_chk102 i_prm_oblgc_chk102(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[102])
);
prm_oblgc_chk103 i_prm_oblgc_chk103(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[103])
);
prm_oblgc_chk104 i_prm_oblgc_chk104(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[104])
);
prm_oblgc_chk105 i_prm_oblgc_chk105(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[105])
);
prm_oblgc_chk106 i_prm_oblgc_chk106(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[106])
);
prm_oblgc_chk107 i_prm_oblgc_chk107(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[107])
);
prm_oblgc_chk108 i_prm_oblgc_chk108(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[108])
);
prm_oblgc_chk109 i_prm_oblgc_chk109(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[109])
);
prm_oblgc_chk110 i_prm_oblgc_chk110(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[110])
);
prm_oblgc_chk111 i_prm_oblgc_chk111(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[111])
);
prm_oblgc_chk112 i_prm_oblgc_chk112(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[112])
);
prm_oblgc_chk113 i_prm_oblgc_chk113(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[113])
);
prm_oblgc_chk114 i_prm_oblgc_chk114(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[114])
);
prm_oblgc_chk115 i_prm_oblgc_chk115(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[115])
);
prm_oblgc_chk116 i_prm_oblgc_chk116(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[116])
);
prm_oblgc_chk117 i_prm_oblgc_chk117(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[117])
);
prm_oblgc_chk118 i_prm_oblgc_chk118(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[118])
);
prm_oblgc_chk119 i_prm_oblgc_chk119(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[119])
);
prm_oblgc_chk120 i_prm_oblgc_chk120(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[120])
);
prm_oblgc_chk121 i_prm_oblgc_chk121(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[121])
);
prm_oblgc_chk122 i_prm_oblgc_chk122(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[122])
);
prm_oblgc_chk123 i_prm_oblgc_chk123(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[123])
);
prm_oblgc_chk124 i_prm_oblgc_chk124(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[124])
);
prm_oblgc_chk125 i_prm_oblgc_chk125(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[125])
);
prm_oblgc_chk126 i_prm_oblgc_chk126(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[126])
);
prm_oblgc_chk127 i_prm_oblgc_chk127(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[127])
);
prm_oblgc_chk128 i_prm_oblgc_chk128(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[128])
);
prm_oblgc_chk129 i_prm_oblgc_chk129(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[129])
);
prm_oblgc_chk130 i_prm_oblgc_chk130(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[130])
);
prm_oblgc_chk131 i_prm_oblgc_chk131(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[131])
);
prm_oblgc_chk132 i_prm_oblgc_chk132(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[132])
);
prm_oblgc_chk133 i_prm_oblgc_chk133(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[133])
);
prm_oblgc_chk134 i_prm_oblgc_chk134(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[134])
);
prm_oblgc_chk135 i_prm_oblgc_chk135(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[135])
);
prm_oblgc_chk136 i_prm_oblgc_chk136(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[136])
);
prm_oblgc_chk137 i_prm_oblgc_chk137(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[137])
);
prm_oblgc_chk138 i_prm_oblgc_chk138(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[138])
);
prm_oblgc_chk139 i_prm_oblgc_chk139(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[139])
);
prm_oblgc_chk140 i_prm_oblgc_chk140(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[140])
);
prm_oblgc_chk141 i_prm_oblgc_chk141(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[141])
);
prm_oblgc_chk142 i_prm_oblgc_chk142(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[142])
);
prm_oblgc_chk143 i_prm_oblgc_chk143(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[143])
);
prm_oblgc_chk144 i_prm_oblgc_chk144(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[144])
);
prm_oblgc_chk145 i_prm_oblgc_chk145(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[145])
);
prm_oblgc_chk146 i_prm_oblgc_chk146(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[146])
);
prm_oblgc_chk147 i_prm_oblgc_chk147(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[147])
);
prm_oblgc_chk148 i_prm_oblgc_chk148(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[148])
);
prm_oblgc_chk149 i_prm_oblgc_chk149(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[149])
);
prm_oblgc_chk150 i_prm_oblgc_chk150(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[150])
);
prm_oblgc_chk151 i_prm_oblgc_chk151(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[151])
);
prm_oblgc_chk152 i_prm_oblgc_chk152(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[152])
);
prm_oblgc_chk153 i_prm_oblgc_chk153(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[153])
);
prm_oblgc_chk154 i_prm_oblgc_chk154(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[154])
);
prm_oblgc_chk155 i_prm_oblgc_chk155(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[155])
);
prm_oblgc_chk156 i_prm_oblgc_chk156(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[156])
);
prm_oblgc_chk157 i_prm_oblgc_chk157(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[157])
);
prm_oblgc_chk158 i_prm_oblgc_chk158(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[158])
);
prm_oblgc_chk159 i_prm_oblgc_chk159(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[159])
);
prm_oblgc_chk160 i_prm_oblgc_chk160(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[160])
);
prm_oblgc_chk161 i_prm_oblgc_chk161(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[161])
);
prm_oblgc_chk162 i_prm_oblgc_chk162(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[162])
);
prm_oblgc_chk163 i_prm_oblgc_chk163(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[163])
);
prm_oblgc_chk164 i_prm_oblgc_chk164(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[164])
);
prm_oblgc_chk165 i_prm_oblgc_chk165(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[165])
);
prm_oblgc_chk166 i_prm_oblgc_chk166(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[166])
);
prm_oblgc_chk167 i_prm_oblgc_chk167(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[167])
);
prm_oblgc_chk168 i_prm_oblgc_chk168(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[168])
);
prm_oblgc_chk169 i_prm_oblgc_chk169(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[169])
);
prm_oblgc_chk170 i_prm_oblgc_chk170(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[170])
);
prm_oblgc_chk171 i_prm_oblgc_chk171(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[171])
);
prm_oblgc_chk172 i_prm_oblgc_chk172(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[172])
);
prm_oblgc_chk173 i_prm_oblgc_chk173(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[173])
);
prm_oblgc_chk174 i_prm_oblgc_chk174(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[174])
);
prm_oblgc_chk175 i_prm_oblgc_chk175(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[175])
);
prm_oblgc_chk176 i_prm_oblgc_chk176(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[176])
);
prm_oblgc_chk177 i_prm_oblgc_chk177(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[177])
);
prm_oblgc_chk178 i_prm_oblgc_chk178(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[178])
);
prm_oblgc_chk179 i_prm_oblgc_chk179(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[179])
);
prm_oblgc_chk180 i_prm_oblgc_chk180(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[180])
);
prm_oblgc_chk181 i_prm_oblgc_chk181(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[181])
);
prm_oblgc_chk182 i_prm_oblgc_chk182(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[182])
);
prm_oblgc_chk183 i_prm_oblgc_chk183(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[183])
);
prm_oblgc_chk184 i_prm_oblgc_chk184(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[184])
);
prm_oblgc_chk185 i_prm_oblgc_chk185(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[185])
);
prm_oblgc_chk186 i_prm_oblgc_chk186(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[186])
);
prm_oblgc_chk187 i_prm_oblgc_chk187(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[187])
);
prm_oblgc_chk188 i_prm_oblgc_chk188(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[188])
);
prm_oblgc_chk189 i_prm_oblgc_chk189(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[189])
);
prm_oblgc_chk190 i_prm_oblgc_chk190(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[190])
);
prm_oblgc_chk191 i_prm_oblgc_chk191(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[191])
);
prm_oblgc_chk192 i_prm_oblgc_chk192(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[192])
);
prm_oblgc_chk193 i_prm_oblgc_chk193(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[193])
);
prm_oblgc_chk194 i_prm_oblgc_chk194(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[194])
);
prm_oblgc_chk195 i_prm_oblgc_chk195(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[195])
);
prm_oblgc_chk196 i_prm_oblgc_chk196(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[196])
);
prm_oblgc_chk197 i_prm_oblgc_chk197(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[197])
);
prm_oblgc_chk198 i_prm_oblgc_chk198(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[198])
);
prm_oblgc_chk199 i_prm_oblgc_chk199(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[199])
);
prm_oblgc_chk200 i_prm_oblgc_chk200(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[200])
);
prm_oblgc_chk201 i_prm_oblgc_chk201(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[201])
);
prm_oblgc_chk202 i_prm_oblgc_chk202(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[202])
);
prm_oblgc_chk203 i_prm_oblgc_chk203(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[203])
);
prm_oblgc_chk204 i_prm_oblgc_chk204(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[204])
);
prm_oblgc_chk205 i_prm_oblgc_chk205(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[205])
);
prm_oblgc_chk206 i_prm_oblgc_chk206(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[206])
);
prm_oblgc_chk207 i_prm_oblgc_chk207(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[207])
);
prm_oblgc_chk208 i_prm_oblgc_chk208(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[208])
);
prm_oblgc_chk209 i_prm_oblgc_chk209(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[209])
);
prm_oblgc_chk210 i_prm_oblgc_chk210(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[210])
);
prm_oblgc_chk211 i_prm_oblgc_chk211(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[211])
);
prm_oblgc_chk212 i_prm_oblgc_chk212(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[212])
);
prm_oblgc_chk213 i_prm_oblgc_chk213(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[213])
);
prm_oblgc_chk214 i_prm_oblgc_chk214(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[214])
);
prm_oblgc_chk215 i_prm_oblgc_chk215(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[215])
);
prm_oblgc_chk216 i_prm_oblgc_chk216(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[216])
);
prm_oblgc_chk217 i_prm_oblgc_chk217(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[217])
);
prm_oblgc_chk218 i_prm_oblgc_chk218(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[218])
);
prm_oblgc_chk219 i_prm_oblgc_chk219(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[219])
);
prm_oblgc_chk220 i_prm_oblgc_chk220(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[220])
);
prm_oblgc_chk221 i_prm_oblgc_chk221(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[221])
);
prm_oblgc_chk222 i_prm_oblgc_chk222(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[222])
);
prm_oblgc_chk223 i_prm_oblgc_chk223(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[223])
);
prm_oblgc_chk224 i_prm_oblgc_chk224(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[224])
);
prm_oblgc_chk225 i_prm_oblgc_chk225(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[225])
);
prm_oblgc_chk226 i_prm_oblgc_chk226(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[226])
);
prm_oblgc_chk227 i_prm_oblgc_chk227(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[227])
);
prm_oblgc_chk228 i_prm_oblgc_chk228(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[228])
);
prm_oblgc_chk229 i_prm_oblgc_chk229(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[229])
);
prm_oblgc_chk230 i_prm_oblgc_chk230(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[230])
);
prm_oblgc_chk231 i_prm_oblgc_chk231(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[231])
);
prm_oblgc_chk232 i_prm_oblgc_chk232(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[232])
);
prm_oblgc_chk233 i_prm_oblgc_chk233(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[233])
);
prm_oblgc_chk234 i_prm_oblgc_chk234(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[234])
);
prm_oblgc_chk235 i_prm_oblgc_chk235(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[235])
);
prm_oblgc_chk236 i_prm_oblgc_chk236(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[236])
);
prm_oblgc_chk237 i_prm_oblgc_chk237(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[237])
);
prm_oblgc_chk238 i_prm_oblgc_chk238(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[238])
);
prm_oblgc_chk239 i_prm_oblgc_chk239(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[239])
);
prm_oblgc_chk240 i_prm_oblgc_chk240(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[240])
);
prm_oblgc_chk241 i_prm_oblgc_chk241(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[241])
);
prm_oblgc_chk242 i_prm_oblgc_chk242(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[242])
);
prm_oblgc_chk243 i_prm_oblgc_chk243(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[243])
);
prm_oblgc_chk244 i_prm_oblgc_chk244(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[244])
);
prm_oblgc_chk245 i_prm_oblgc_chk245(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[245])
);
prm_oblgc_chk246 i_prm_oblgc_chk246(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[246])
);
prm_oblgc_chk247 i_prm_oblgc_chk247(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[247])
);
prm_oblgc_chk248 i_prm_oblgc_chk248(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[248])
);
prm_oblgc_chk249 i_prm_oblgc_chk249(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[249])
);
prm_oblgc_chk250 i_prm_oblgc_chk250(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[250])
);
prm_oblgc_chk251 i_prm_oblgc_chk251(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[251])
);
prm_oblgc_chk252 i_prm_oblgc_chk252(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[252])
);
prm_oblgc_chk253 i_prm_oblgc_chk253(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[253])
);
prm_oblgc_chk254 i_prm_oblgc_chk254(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[254])
);
prm_oblgc_chk255 i_prm_oblgc_chk255(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[255])
);
prm_oblgc_chk256 i_prm_oblgc_chk256(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[256])
);
prm_oblgc_chk257 i_prm_oblgc_chk257(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[257])
);
prm_oblgc_chk258 i_prm_oblgc_chk258(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[258])
);
prm_oblgc_chk259 i_prm_oblgc_chk259(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[259])
);
prm_oblgc_chk260 i_prm_oblgc_chk260(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[260])
);
prm_oblgc_chk261 i_prm_oblgc_chk261(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[261])
);
prm_oblgc_chk262 i_prm_oblgc_chk262(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[262])
);
prm_oblgc_chk263 i_prm_oblgc_chk263(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[263])
);
prm_oblgc_chk264 i_prm_oblgc_chk264(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[264])
);
prm_oblgc_chk265 i_prm_oblgc_chk265(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[265])
);
prm_oblgc_chk266 i_prm_oblgc_chk266(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[266])
);
prm_oblgc_chk267 i_prm_oblgc_chk267(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[267])
);
prm_oblgc_chk268 i_prm_oblgc_chk268(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[268])
);
prm_oblgc_chk269 i_prm_oblgc_chk269(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[269])
);
prm_oblgc_chk270 i_prm_oblgc_chk270(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[270])
);
prm_oblgc_chk271 i_prm_oblgc_chk271(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[271])
);
prm_oblgc_chk272 i_prm_oblgc_chk272(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[272])
);
prm_oblgc_chk273 i_prm_oblgc_chk273(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[273])
);
prm_oblgc_chk274 i_prm_oblgc_chk274(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[274])
);
prm_oblgc_chk275 i_prm_oblgc_chk275(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[275])
);
prm_oblgc_chk276 i_prm_oblgc_chk276(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[276])
);
prm_oblgc_chk277 i_prm_oblgc_chk277(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[277])
);
prm_oblgc_chk278 i_prm_oblgc_chk278(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[278])
);
prm_oblgc_chk279 i_prm_oblgc_chk279(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[279])
);
prm_oblgc_chk280 i_prm_oblgc_chk280(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[280])
);
prm_oblgc_chk281 i_prm_oblgc_chk281(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[281])
);
prm_oblgc_chk282 i_prm_oblgc_chk282(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[282])
);
prm_oblgc_chk283 i_prm_oblgc_chk283(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[283])
);
prm_oblgc_chk284 i_prm_oblgc_chk284(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[284])
);
prm_oblgc_chk285 i_prm_oblgc_chk285(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[285])
);
prm_oblgc_chk286 i_prm_oblgc_chk286(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[286])
);
prm_oblgc_chk287 i_prm_oblgc_chk287(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[287])
);
prm_oblgc_chk288 i_prm_oblgc_chk288(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[288])
);
prm_oblgc_chk289 i_prm_oblgc_chk289(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[289])
);
prm_oblgc_chk290 i_prm_oblgc_chk290(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[290])
);
prm_oblgc_chk291 i_prm_oblgc_chk291(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[291])
);
prm_oblgc_chk292 i_prm_oblgc_chk292(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[292])
);
prm_oblgc_chk293 i_prm_oblgc_chk293(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[293])
);
prm_oblgc_chk294 i_prm_oblgc_chk294(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[294])
);
prm_oblgc_chk295 i_prm_oblgc_chk295(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[295])
);
prm_oblgc_chk296 i_prm_oblgc_chk296(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[296])
);
prm_oblgc_chk297 i_prm_oblgc_chk297(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[297])
);
prm_oblgc_chk298 i_prm_oblgc_chk298(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[298])
);
prm_oblgc_chk299 i_prm_oblgc_chk299(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[299])
);
prm_oblgc_chk300 i_prm_oblgc_chk300(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[300])
);
prm_oblgc_chk301 i_prm_oblgc_chk301(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[301])
);
prm_oblgc_chk302 i_prm_oblgc_chk302(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[302])
);
prm_oblgc_chk303 i_prm_oblgc_chk303(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[303])
);
prm_oblgc_chk304 i_prm_oblgc_chk304(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[304])
);
prm_oblgc_chk305 i_prm_oblgc_chk305(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[305])
);
prm_oblgc_chk306 i_prm_oblgc_chk306(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[306])
);
prm_oblgc_chk307 i_prm_oblgc_chk307(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[307])
);
prm_oblgc_chk308 i_prm_oblgc_chk308(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[308])
);
prm_oblgc_chk309 i_prm_oblgc_chk309(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[309])
);
prm_oblgc_chk310 i_prm_oblgc_chk310(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[310])
);
prm_oblgc_chk311 i_prm_oblgc_chk311(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[311])
);
prm_oblgc_chk312 i_prm_oblgc_chk312(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[312])
);
prm_oblgc_chk313 i_prm_oblgc_chk313(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[313])
);
prm_oblgc_chk314 i_prm_oblgc_chk314(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[314])
);
prm_oblgc_chk315 i_prm_oblgc_chk315(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[315])
);
prm_oblgc_chk316 i_prm_oblgc_chk316(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[316])
);
prm_oblgc_chk317 i_prm_oblgc_chk317(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[317])
);
prm_oblgc_chk318 i_prm_oblgc_chk318(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[318])
);
prm_oblgc_chk319 i_prm_oblgc_chk319(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[319])
);
prm_oblgc_chk320 i_prm_oblgc_chk320(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[320])
);
prm_oblgc_chk321 i_prm_oblgc_chk321(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[321])
);
prm_oblgc_chk322 i_prm_oblgc_chk322(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[322])
);
prm_oblgc_chk323 i_prm_oblgc_chk323(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[323])
);
prm_oblgc_chk324 i_prm_oblgc_chk324(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[324])
);
prm_oblgc_chk325 i_prm_oblgc_chk325(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[325])
);
prm_oblgc_chk326 i_prm_oblgc_chk326(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[326])
);
prm_oblgc_chk327 i_prm_oblgc_chk327(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[327])
);
prm_oblgc_chk328 i_prm_oblgc_chk328(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[328])
);
prm_oblgc_chk329 i_prm_oblgc_chk329(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[329])
);
prm_oblgc_chk330 i_prm_oblgc_chk330(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[330])
);
prm_oblgc_chk331 i_prm_oblgc_chk331(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[331])
);
prm_oblgc_chk332 i_prm_oblgc_chk332(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[332])
);
prm_oblgc_chk333 i_prm_oblgc_chk333(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[333])
);
prm_oblgc_chk334 i_prm_oblgc_chk334(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[334])
);
prm_oblgc_chk335 i_prm_oblgc_chk335(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[335])
);
prm_oblgc_chk336 i_prm_oblgc_chk336(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[336])
);
prm_oblgc_chk337 i_prm_oblgc_chk337(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[337])
);
prm_oblgc_chk338 i_prm_oblgc_chk338(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[338])
);
prm_oblgc_chk339 i_prm_oblgc_chk339(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[339])
);
prm_oblgc_chk340 i_prm_oblgc_chk340(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[340])
);
prm_oblgc_chk341 i_prm_oblgc_chk341(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[341])
);
prm_oblgc_chk342 i_prm_oblgc_chk342(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[342])
);
prm_oblgc_chk343 i_prm_oblgc_chk343(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[343])
);
prm_oblgc_chk344 i_prm_oblgc_chk344(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[344])
);
prm_oblgc_chk345 i_prm_oblgc_chk345(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[345])
);
prm_oblgc_chk346 i_prm_oblgc_chk346(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[346])
);
prm_oblgc_chk347 i_prm_oblgc_chk347(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[347])
);
prm_oblgc_chk348 i_prm_oblgc_chk348(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[348])
);
prm_oblgc_chk349 i_prm_oblgc_chk349(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[349])
);
prm_oblgc_chk350 i_prm_oblgc_chk350(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[350])
);
prm_oblgc_chk351 i_prm_oblgc_chk351(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[351])
);
prm_oblgc_chk352 i_prm_oblgc_chk352(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[352])
);
prm_oblgc_chk353 i_prm_oblgc_chk353(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[353])
);
prm_oblgc_chk354 i_prm_oblgc_chk354(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[354])
);
prm_oblgc_chk355 i_prm_oblgc_chk355(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[355])
);
prm_oblgc_chk356 i_prm_oblgc_chk356(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[356])
);
prm_oblgc_chk357 i_prm_oblgc_chk357(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[357])
);
prm_oblgc_chk358 i_prm_oblgc_chk358(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[358])
);
prm_oblgc_chk359 i_prm_oblgc_chk359(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[359])
);
prm_oblgc_chk360 i_prm_oblgc_chk360(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[360])
);
prm_oblgc_chk361 i_prm_oblgc_chk361(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[361])
);
prm_oblgc_chk362 i_prm_oblgc_chk362(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[362])
);
prm_oblgc_chk363 i_prm_oblgc_chk363(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[363])
);
prm_oblgc_chk364 i_prm_oblgc_chk364(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[364])
);
prm_oblgc_chk365 i_prm_oblgc_chk365(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[365])
);
prm_oblgc_chk366 i_prm_oblgc_chk366(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[366])
);
prm_oblgc_chk367 i_prm_oblgc_chk367(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[367])
);
prm_oblgc_chk368 i_prm_oblgc_chk368(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[368])
);
prm_oblgc_chk369 i_prm_oblgc_chk369(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[369])
);
prm_oblgc_chk370 i_prm_oblgc_chk370(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[370])
);
prm_oblgc_chk371 i_prm_oblgc_chk371(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[371])
);
prm_oblgc_chk372 i_prm_oblgc_chk372(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[372])
);
prm_oblgc_chk373 i_prm_oblgc_chk373(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[373])
);
prm_oblgc_chk374 i_prm_oblgc_chk374(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[374])
);
prm_oblgc_chk375 i_prm_oblgc_chk375(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[375])
);
prm_oblgc_chk376 i_prm_oblgc_chk376(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[376])
);
prm_oblgc_chk377 i_prm_oblgc_chk377(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[377])
);
prm_oblgc_chk378 i_prm_oblgc_chk378(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[378])
);
prm_oblgc_chk379 i_prm_oblgc_chk379(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[379])
);
prm_oblgc_chk380 i_prm_oblgc_chk380(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[380])
);
prm_oblgc_chk381 i_prm_oblgc_chk381(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[381])
);
prm_oblgc_chk382 i_prm_oblgc_chk382(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[382])
);
prm_oblgc_chk383 i_prm_oblgc_chk383(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[383])
);
prm_oblgc_chk384 i_prm_oblgc_chk384(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[384])
);
prm_oblgc_chk385 i_prm_oblgc_chk385(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[385])
);
prm_oblgc_chk386 i_prm_oblgc_chk386(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[386])
);
prm_oblgc_chk387 i_prm_oblgc_chk387(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[387])
);
prm_oblgc_chk388 i_prm_oblgc_chk388(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[388])
);
prm_oblgc_chk389 i_prm_oblgc_chk389(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[389])
);
prm_oblgc_chk390 i_prm_oblgc_chk390(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[390])
);
prm_oblgc_chk391 i_prm_oblgc_chk391(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[391])
);
prm_oblgc_chk392 i_prm_oblgc_chk392(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[392])
);
prm_oblgc_chk393 i_prm_oblgc_chk393(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[393])
);
prm_oblgc_chk394 i_prm_oblgc_chk394(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[394])
);
prm_oblgc_chk395 i_prm_oblgc_chk395(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[395])
);
prm_oblgc_chk396 i_prm_oblgc_chk396(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[396])
);
prm_oblgc_chk397 i_prm_oblgc_chk397(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[397])
);
prm_oblgc_chk398 i_prm_oblgc_chk398(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[398])
);
prm_oblgc_chk399 i_prm_oblgc_chk399(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[399])
);
prm_oblgc_chk400 i_prm_oblgc_chk400(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[400])
);
prm_oblgc_chk401 i_prm_oblgc_chk401(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[401])
);
prm_oblgc_chk402 i_prm_oblgc_chk402(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[402])
);
prm_oblgc_chk403 i_prm_oblgc_chk403(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[403])
);
prm_oblgc_chk404 i_prm_oblgc_chk404(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[404])
);
prm_oblgc_chk405 i_prm_oblgc_chk405(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[405])
);
prm_oblgc_chk406 i_prm_oblgc_chk406(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[406])
);
prm_oblgc_chk407 i_prm_oblgc_chk407(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[407])
);
prm_oblgc_chk408 i_prm_oblgc_chk408(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[408])
);
prm_oblgc_chk409 i_prm_oblgc_chk409(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[409])
);
prm_oblgc_chk410 i_prm_oblgc_chk410(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[410])
);
prm_oblgc_chk411 i_prm_oblgc_chk411(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[411])
);
prm_oblgc_chk412 i_prm_oblgc_chk412(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[412])
);
prm_oblgc_chk413 i_prm_oblgc_chk413(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[413])
);
prm_oblgc_chk414 i_prm_oblgc_chk414(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[414])
);
prm_oblgc_chk415 i_prm_oblgc_chk415(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[415])
);
prm_oblgc_chk416 i_prm_oblgc_chk416(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[416])
);
prm_oblgc_chk417 i_prm_oblgc_chk417(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[417])
);
prm_oblgc_chk418 i_prm_oblgc_chk418(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[418])
);
prm_oblgc_chk419 i_prm_oblgc_chk419(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[419])
);
prm_oblgc_chk420 i_prm_oblgc_chk420(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[420])
);
prm_oblgc_chk421 i_prm_oblgc_chk421(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[421])
);
prm_oblgc_chk422 i_prm_oblgc_chk422(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[422])
);
prm_oblgc_chk423 i_prm_oblgc_chk423(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[423])
);
prm_oblgc_chk424 i_prm_oblgc_chk424(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[424])
);
prm_oblgc_chk425 i_prm_oblgc_chk425(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[425])
);
prm_oblgc_chk426 i_prm_oblgc_chk426(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[426])
);
prm_oblgc_chk427 i_prm_oblgc_chk427(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[427])
);
prm_oblgc_chk428 i_prm_oblgc_chk428(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[428])
);
prm_oblgc_chk429 i_prm_oblgc_chk429(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[429])
);
prm_oblgc_chk430 i_prm_oblgc_chk430(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[430])
);
prm_oblgc_chk431 i_prm_oblgc_chk431(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[431])
);
prm_oblgc_chk432 i_prm_oblgc_chk432(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[432])
);
prm_oblgc_chk433 i_prm_oblgc_chk433(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[433])
);
prm_oblgc_chk434 i_prm_oblgc_chk434(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[434])
);
prm_oblgc_chk435 i_prm_oblgc_chk435(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[435])
);
prm_oblgc_chk436 i_prm_oblgc_chk436(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[436])
);
prm_oblgc_chk437 i_prm_oblgc_chk437(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[437])
);
prm_oblgc_chk438 i_prm_oblgc_chk438(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[438])
);
prm_oblgc_chk439 i_prm_oblgc_chk439(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[439])
);
prm_oblgc_chk440 i_prm_oblgc_chk440(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[440])
);
prm_oblgc_chk441 i_prm_oblgc_chk441(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[441])
);
prm_oblgc_chk442 i_prm_oblgc_chk442(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[442])
);
prm_oblgc_chk443 i_prm_oblgc_chk443(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[443])
);
prm_oblgc_chk444 i_prm_oblgc_chk444(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[444])
);
prm_oblgc_chk445 i_prm_oblgc_chk445(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[445])
);
prm_oblgc_chk446 i_prm_oblgc_chk446(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[446])
);
prm_oblgc_chk447 i_prm_oblgc_chk447(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[447])
);
prm_oblgc_chk448 i_prm_oblgc_chk448(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[448])
);
prm_oblgc_chk449 i_prm_oblgc_chk449(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[449])
);
prm_oblgc_chk450 i_prm_oblgc_chk450(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[450])
);
prm_oblgc_chk451 i_prm_oblgc_chk451(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[451])
);
prm_oblgc_chk452 i_prm_oblgc_chk452(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[452])
);
prm_oblgc_chk453 i_prm_oblgc_chk453(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[453])
);
prm_oblgc_chk454 i_prm_oblgc_chk454(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[454])
);
prm_oblgc_chk455 i_prm_oblgc_chk455(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[455])
);
prm_oblgc_chk456 i_prm_oblgc_chk456(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[456])
);
prm_oblgc_chk457 i_prm_oblgc_chk457(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[457])
);
prm_oblgc_chk458 i_prm_oblgc_chk458(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[458])
);
prm_oblgc_chk459 i_prm_oblgc_chk459(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[459])
);
prm_oblgc_chk460 i_prm_oblgc_chk460(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[460])
);
prm_oblgc_chk461 i_prm_oblgc_chk461(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[461])
);
prm_oblgc_chk462 i_prm_oblgc_chk462(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[462])
);
prm_oblgc_chk463 i_prm_oblgc_chk463(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[463])
);
prm_oblgc_chk464 i_prm_oblgc_chk464(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[464])
);
prm_oblgc_chk465 i_prm_oblgc_chk465(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[465])
);
prm_oblgc_chk466 i_prm_oblgc_chk466(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[466])
);
prm_oblgc_chk467 i_prm_oblgc_chk467(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[467])
);
prm_oblgc_chk468 i_prm_oblgc_chk468(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[468])
);
prm_oblgc_chk469 i_prm_oblgc_chk469(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[469])
);
prm_oblgc_chk470 i_prm_oblgc_chk470(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[470])
);
prm_oblgc_chk471 i_prm_oblgc_chk471(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[471])
);
prm_oblgc_chk472 i_prm_oblgc_chk472(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[472])
);
prm_oblgc_chk473 i_prm_oblgc_chk473(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[473])
);
prm_oblgc_chk474 i_prm_oblgc_chk474(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[474])
);
prm_oblgc_chk475 i_prm_oblgc_chk475(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[475])
);
prm_oblgc_chk476 i_prm_oblgc_chk476(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[476])
);
prm_oblgc_chk477 i_prm_oblgc_chk477(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[477])
);
prm_oblgc_chk478 i_prm_oblgc_chk478(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[478])
);
prm_oblgc_chk479 i_prm_oblgc_chk479(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[479])
);
prm_oblgc_chk480 i_prm_oblgc_chk480(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[480])
);
prm_oblgc_chk481 i_prm_oblgc_chk481(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[481])
);
prm_oblgc_chk482 i_prm_oblgc_chk482(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[482])
);
prm_oblgc_chk483 i_prm_oblgc_chk483(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[483])
);
prm_oblgc_chk484 i_prm_oblgc_chk484(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[484])
);
prm_oblgc_chk485 i_prm_oblgc_chk485(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[485])
);
prm_oblgc_chk486 i_prm_oblgc_chk486(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[486])
);
prm_oblgc_chk487 i_prm_oblgc_chk487(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[487])
);
prm_oblgc_chk488 i_prm_oblgc_chk488(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[488])
);
prm_oblgc_chk489 i_prm_oblgc_chk489(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[489])
);
prm_oblgc_chk490 i_prm_oblgc_chk490(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[490])
);
prm_oblgc_chk491 i_prm_oblgc_chk491(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[491])
);
prm_oblgc_chk492 i_prm_oblgc_chk492(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[492])
);
prm_oblgc_chk493 i_prm_oblgc_chk493(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[493])
);
prm_oblgc_chk494 i_prm_oblgc_chk494(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[494])
);
prm_oblgc_chk495 i_prm_oblgc_chk495(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[495])
);
prm_oblgc_chk496 i_prm_oblgc_chk496(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[496])
);
prm_oblgc_chk497 i_prm_oblgc_chk497(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[497])
);
prm_oblgc_chk498 i_prm_oblgc_chk498(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[498])
);
prm_oblgc_chk499 i_prm_oblgc_chk499(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[499])
);
prm_oblgc_chk500 i_prm_oblgc_chk500(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[500])
);
prm_oblgc_chk501 i_prm_oblgc_chk501(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[501])
);
prm_oblgc_chk502 i_prm_oblgc_chk502(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[502])
);
prm_oblgc_chk503 i_prm_oblgc_chk503(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[503])
);
prm_oblgc_chk504 i_prm_oblgc_chk504(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[504])
);
prm_oblgc_chk505 i_prm_oblgc_chk505(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[505])
);
prm_oblgc_chk506 i_prm_oblgc_chk506(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[506])
);
prm_oblgc_chk507 i_prm_oblgc_chk507(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[507])
);
prm_oblgc_chk508 i_prm_oblgc_chk508(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[508])
);
prm_oblgc_chk509 i_prm_oblgc_chk509(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[509])
);
prm_oblgc_chk510 i_prm_oblgc_chk510(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[510])
);
prm_oblgc_chk511 i_prm_oblgc_chk511(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[511])
);
prm_oblgc_chk512 i_prm_oblgc_chk512(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[512])
);
prm_oblgc_chk513 i_prm_oblgc_chk513(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[513])
);
prm_oblgc_chk514 i_prm_oblgc_chk514(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[514])
);
prm_oblgc_chk515 i_prm_oblgc_chk515(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[515])
);
prm_oblgc_chk516 i_prm_oblgc_chk516(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[516])
);
prm_oblgc_chk517 i_prm_oblgc_chk517(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[517])
);
prm_oblgc_chk518 i_prm_oblgc_chk518(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[518])
);
prm_oblgc_chk519 i_prm_oblgc_chk519(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[519])
);
prm_oblgc_chk520 i_prm_oblgc_chk520(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[520])
);
prm_oblgc_chk521 i_prm_oblgc_chk521(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[521])
);
prm_oblgc_chk522 i_prm_oblgc_chk522(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[522])
);
prm_oblgc_chk523 i_prm_oblgc_chk523(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[523])
);
prm_oblgc_chk524 i_prm_oblgc_chk524(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[524])
);
prm_oblgc_chk525 i_prm_oblgc_chk525(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[525])
);
prm_oblgc_chk526 i_prm_oblgc_chk526(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[526])
);
prm_oblgc_chk527 i_prm_oblgc_chk527(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[527])
);
prm_oblgc_chk528 i_prm_oblgc_chk528(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[528])
);
prm_oblgc_chk529 i_prm_oblgc_chk529(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[529])
);
prm_oblgc_chk530 i_prm_oblgc_chk530(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[530])
);
prm_oblgc_chk531 i_prm_oblgc_chk531(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[531])
);
prm_oblgc_chk532 i_prm_oblgc_chk532(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[532])
);
prm_oblgc_chk533 i_prm_oblgc_chk533(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[533])
);
prm_oblgc_chk534 i_prm_oblgc_chk534(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[534])
);
prm_oblgc_chk535 i_prm_oblgc_chk535(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[535])
);
prm_oblgc_chk536 i_prm_oblgc_chk536(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[536])
);
prm_oblgc_chk537 i_prm_oblgc_chk537(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[537])
);
prm_oblgc_chk538 i_prm_oblgc_chk538(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[538])
);
prm_oblgc_chk539 i_prm_oblgc_chk539(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[539])
);
prm_oblgc_chk540 i_prm_oblgc_chk540(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[540])
);
prm_oblgc_chk541 i_prm_oblgc_chk541(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[541])
);
prm_oblgc_chk542 i_prm_oblgc_chk542(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[542])
);
prm_oblgc_chk543 i_prm_oblgc_chk543(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[543])
);
prm_oblgc_chk544 i_prm_oblgc_chk544(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[544])
);
prm_oblgc_chk545 i_prm_oblgc_chk545(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[545])
);
prm_oblgc_chk546 i_prm_oblgc_chk546(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[546])
);
prm_oblgc_chk547 i_prm_oblgc_chk547(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[547])
);
prm_oblgc_chk548 i_prm_oblgc_chk548(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[548])
);
prm_oblgc_chk549 i_prm_oblgc_chk549(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[549])
);
prm_oblgc_chk550 i_prm_oblgc_chk550(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[550])
);
prm_oblgc_chk551 i_prm_oblgc_chk551(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[551])
);
prm_oblgc_chk552 i_prm_oblgc_chk552(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[552])
);
prm_oblgc_chk553 i_prm_oblgc_chk553(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[553])
);
prm_oblgc_chk554 i_prm_oblgc_chk554(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[554])
);
prm_oblgc_chk555 i_prm_oblgc_chk555(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[555])
);
prm_oblgc_chk556 i_prm_oblgc_chk556(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[556])
);
prm_oblgc_chk557 i_prm_oblgc_chk557(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[557])
);
prm_oblgc_chk558 i_prm_oblgc_chk558(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[558])
);
prm_oblgc_chk559 i_prm_oblgc_chk559(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[559])
);
prm_oblgc_chk560 i_prm_oblgc_chk560(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[560])
);
prm_oblgc_chk561 i_prm_oblgc_chk561(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[561])
);
prm_oblgc_chk562 i_prm_oblgc_chk562(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[562])
);
prm_oblgc_chk563 i_prm_oblgc_chk563(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[563])
);
prm_oblgc_chk564 i_prm_oblgc_chk564(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[564])
);
prm_oblgc_chk565 i_prm_oblgc_chk565(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[565])
);
prm_oblgc_chk566 i_prm_oblgc_chk566(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[566])
);
prm_oblgc_chk567 i_prm_oblgc_chk567(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[567])
);
prm_oblgc_chk568 i_prm_oblgc_chk568(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[568])
);
prm_oblgc_chk569 i_prm_oblgc_chk569(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[569])
);
prm_oblgc_chk570 i_prm_oblgc_chk570(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[570])
);
prm_oblgc_chk571 i_prm_oblgc_chk571(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[571])
);
prm_oblgc_chk572 i_prm_oblgc_chk572(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[572])
);
prm_oblgc_chk573 i_prm_oblgc_chk573(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[573])
);
prm_oblgc_chk574 i_prm_oblgc_chk574(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[574])
);
prm_oblgc_chk575 i_prm_oblgc_chk575(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[575])
);
prm_oblgc_chk576 i_prm_oblgc_chk576(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[576])
);
prm_oblgc_chk577 i_prm_oblgc_chk577(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[577])
);
prm_oblgc_chk578 i_prm_oblgc_chk578(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[578])
);
prm_oblgc_chk579 i_prm_oblgc_chk579(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[579])
);
prm_oblgc_chk580 i_prm_oblgc_chk580(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[580])
);
prm_oblgc_chk581 i_prm_oblgc_chk581(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[581])
);
prm_oblgc_chk582 i_prm_oblgc_chk582(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[582])
);
prm_oblgc_chk583 i_prm_oblgc_chk583(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[583])
);
prm_oblgc_chk584 i_prm_oblgc_chk584(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[584])
);
prm_oblgc_chk585 i_prm_oblgc_chk585(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[585])
);
prm_oblgc_chk586 i_prm_oblgc_chk586(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[586])
);
prm_oblgc_chk587 i_prm_oblgc_chk587(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[587])
);
prm_oblgc_chk588 i_prm_oblgc_chk588(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[588])
);
prm_oblgc_chk589 i_prm_oblgc_chk589(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[589])
);
prm_oblgc_chk590 i_prm_oblgc_chk590(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[590])
);
prm_oblgc_chk591 i_prm_oblgc_chk591(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[591])
);
prm_oblgc_chk592 i_prm_oblgc_chk592(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[592])
);
prm_oblgc_chk593 i_prm_oblgc_chk593(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[593])
);
prm_oblgc_chk594 i_prm_oblgc_chk594(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[594])
);
prm_oblgc_chk595 i_prm_oblgc_chk595(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[595])
);
prm_oblgc_chk596 i_prm_oblgc_chk596(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[596])
);
prm_oblgc_chk597 i_prm_oblgc_chk597(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[597])
);
prm_oblgc_chk598 i_prm_oblgc_chk598(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[598])
);
prm_oblgc_chk599 i_prm_oblgc_chk599(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[599])
);
prm_oblgc_chk600 i_prm_oblgc_chk600(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[600])
);
prm_oblgc_chk601 i_prm_oblgc_chk601(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[601])
);
prm_oblgc_chk602 i_prm_oblgc_chk602(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[602])
);
prm_oblgc_chk603 i_prm_oblgc_chk603(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[603])
);
prm_oblgc_chk604 i_prm_oblgc_chk604(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[604])
);
prm_oblgc_chk605 i_prm_oblgc_chk605(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[605])
);
prm_oblgc_chk606 i_prm_oblgc_chk606(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[606])
);
prm_oblgc_chk607 i_prm_oblgc_chk607(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[607])
);
prm_oblgc_chk608 i_prm_oblgc_chk608(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[608])
);
prm_oblgc_chk609 i_prm_oblgc_chk609(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[609])
);
prm_oblgc_chk610 i_prm_oblgc_chk610(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[610])
);
prm_oblgc_chk611 i_prm_oblgc_chk611(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[611])
);
prm_oblgc_chk612 i_prm_oblgc_chk612(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[612])
);
prm_oblgc_chk613 i_prm_oblgc_chk613(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[613])
);
prm_oblgc_chk614 i_prm_oblgc_chk614(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[614])
);
prm_oblgc_chk615 i_prm_oblgc_chk615(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[615])
);
prm_oblgc_chk616 i_prm_oblgc_chk616(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[616])
);
prm_oblgc_chk617 i_prm_oblgc_chk617(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[617])
);
prm_oblgc_chk618 i_prm_oblgc_chk618(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[618])
);
prm_oblgc_chk619 i_prm_oblgc_chk619(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[619])
);
prm_oblgc_chk620 i_prm_oblgc_chk620(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[620])
);
prm_oblgc_chk621 i_prm_oblgc_chk621(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[621])
);
prm_oblgc_chk622 i_prm_oblgc_chk622(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[622])
);
prm_oblgc_chk623 i_prm_oblgc_chk623(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[623])
);
prm_oblgc_chk624 i_prm_oblgc_chk624(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[624])
);
prm_oblgc_chk625 i_prm_oblgc_chk625(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[625])
);
prm_oblgc_chk626 i_prm_oblgc_chk626(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[626])
);
prm_oblgc_chk627 i_prm_oblgc_chk627(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[627])
);
prm_oblgc_chk628 i_prm_oblgc_chk628(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[628])
);
prm_oblgc_chk629 i_prm_oblgc_chk629(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[629])
);
prm_oblgc_chk630 i_prm_oblgc_chk630(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[630])
);
prm_oblgc_chk631 i_prm_oblgc_chk631(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[631])
);
prm_oblgc_chk632 i_prm_oblgc_chk632(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[632])
);
prm_oblgc_chk633 i_prm_oblgc_chk633(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[633])
);
prm_oblgc_chk634 i_prm_oblgc_chk634(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[634])
);
prm_oblgc_chk635 i_prm_oblgc_chk635(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[635])
);
prm_oblgc_chk636 i_prm_oblgc_chk636(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[636])
);
prm_oblgc_chk637 i_prm_oblgc_chk637(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[637])
);
prm_oblgc_chk638 i_prm_oblgc_chk638(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[638])
);
prm_oblgc_chk639 i_prm_oblgc_chk639(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[639])
);
prm_oblgc_chk640 i_prm_oblgc_chk640(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[640])
);
prm_oblgc_chk641 i_prm_oblgc_chk641(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[641])
);
prm_oblgc_chk642 i_prm_oblgc_chk642(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[642])
);
prm_oblgc_chk643 i_prm_oblgc_chk643(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[643])
);
prm_oblgc_chk644 i_prm_oblgc_chk644(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[644])
);
prm_oblgc_chk645 i_prm_oblgc_chk645(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[645])
);
prm_oblgc_chk646 i_prm_oblgc_chk646(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[646])
);
prm_oblgc_chk647 i_prm_oblgc_chk647(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[647])
);
prm_oblgc_chk648 i_prm_oblgc_chk648(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[648])
);
prm_oblgc_chk649 i_prm_oblgc_chk649(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[649])
);
prm_oblgc_chk650 i_prm_oblgc_chk650(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[650])
);
prm_oblgc_chk651 i_prm_oblgc_chk651(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[651])
);
prm_oblgc_chk652 i_prm_oblgc_chk652(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[652])
);
prm_oblgc_chk653 i_prm_oblgc_chk653(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[653])
);
prm_oblgc_chk654 i_prm_oblgc_chk654(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[654])
);
prm_oblgc_chk655 i_prm_oblgc_chk655(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[655])
);
prm_oblgc_chk656 i_prm_oblgc_chk656(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[656])
);
prm_oblgc_chk657 i_prm_oblgc_chk657(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[657])
);
prm_oblgc_chk658 i_prm_oblgc_chk658(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[658])
);
prm_oblgc_chk659 i_prm_oblgc_chk659(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[659])
);
prm_oblgc_chk660 i_prm_oblgc_chk660(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[660])
);
prm_oblgc_chk661 i_prm_oblgc_chk661(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[661])
);
prm_oblgc_chk662 i_prm_oblgc_chk662(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[662])
);
prm_oblgc_chk663 i_prm_oblgc_chk663(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[663])
);
prm_oblgc_chk664 i_prm_oblgc_chk664(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[664])
);
prm_oblgc_chk665 i_prm_oblgc_chk665(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[665])
);
prm_oblgc_chk666 i_prm_oblgc_chk666(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[666])
);
prm_oblgc_chk667 i_prm_oblgc_chk667(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[667])
);
prm_oblgc_chk668 i_prm_oblgc_chk668(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[668])
);
prm_oblgc_chk669 i_prm_oblgc_chk669(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[669])
);
prm_oblgc_chk670 i_prm_oblgc_chk670(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[670])
);
prm_oblgc_chk671 i_prm_oblgc_chk671(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[671])
);
prm_oblgc_chk672 i_prm_oblgc_chk672(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[672])
);
prm_oblgc_chk673 i_prm_oblgc_chk673(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[673])
);
prm_oblgc_chk674 i_prm_oblgc_chk674(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[674])
);
prm_oblgc_chk675 i_prm_oblgc_chk675(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[675])
);
prm_oblgc_chk676 i_prm_oblgc_chk676(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[676])
);
prm_oblgc_chk677 i_prm_oblgc_chk677(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[677])
);
prm_oblgc_chk678 i_prm_oblgc_chk678(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[678])
);
prm_oblgc_chk679 i_prm_oblgc_chk679(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[679])
);
prm_oblgc_chk680 i_prm_oblgc_chk680(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[680])
);
prm_oblgc_chk681 i_prm_oblgc_chk681(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[681])
);
prm_oblgc_chk682 i_prm_oblgc_chk682(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[682])
);
prm_oblgc_chk683 i_prm_oblgc_chk683(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[683])
);
prm_oblgc_chk684 i_prm_oblgc_chk684(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[684])
);
prm_oblgc_chk685 i_prm_oblgc_chk685(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[685])
);
prm_oblgc_chk686 i_prm_oblgc_chk686(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[686])
);
prm_oblgc_chk687 i_prm_oblgc_chk687(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[687])
);
prm_oblgc_chk688 i_prm_oblgc_chk688(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[688])
);
prm_oblgc_chk689 i_prm_oblgc_chk689(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[689])
);
prm_oblgc_chk690 i_prm_oblgc_chk690(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[690])
);
prm_oblgc_chk691 i_prm_oblgc_chk691(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[691])
);
prm_oblgc_chk692 i_prm_oblgc_chk692(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[692])
);
prm_oblgc_chk693 i_prm_oblgc_chk693(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[693])
);
prm_oblgc_chk694 i_prm_oblgc_chk694(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[694])
);
prm_oblgc_chk695 i_prm_oblgc_chk695(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[695])
);
prm_oblgc_chk696 i_prm_oblgc_chk696(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[696])
);
prm_oblgc_chk697 i_prm_oblgc_chk697(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[697])
);
prm_oblgc_chk698 i_prm_oblgc_chk698(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[698])
);
prm_oblgc_chk699 i_prm_oblgc_chk699(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[699])
);
prm_oblgc_chk700 i_prm_oblgc_chk700(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[700])
);
prm_oblgc_chk701 i_prm_oblgc_chk701(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[701])
);
prm_oblgc_chk702 i_prm_oblgc_chk702(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[702])
);
prm_oblgc_chk703 i_prm_oblgc_chk703(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[703])
);
prm_oblgc_chk704 i_prm_oblgc_chk704(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[704])
);
prm_oblgc_chk705 i_prm_oblgc_chk705(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[705])
);
prm_oblgc_chk706 i_prm_oblgc_chk706(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[706])
);
prm_oblgc_chk707 i_prm_oblgc_chk707(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[707])
);
prm_oblgc_chk708 i_prm_oblgc_chk708(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[708])
);
prm_oblgc_chk709 i_prm_oblgc_chk709(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[709])
);
prm_oblgc_chk710 i_prm_oblgc_chk710(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[710])
);
prm_oblgc_chk711 i_prm_oblgc_chk711(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[711])
);
prm_oblgc_chk712 i_prm_oblgc_chk712(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[712])
);
prm_oblgc_chk713 i_prm_oblgc_chk713(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[713])
);
prm_oblgc_chk714 i_prm_oblgc_chk714(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[714])
);
prm_oblgc_chk715 i_prm_oblgc_chk715(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[715])
);
prm_oblgc_chk716 i_prm_oblgc_chk716(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[716])
);
prm_oblgc_chk717 i_prm_oblgc_chk717(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[717])
);
prm_oblgc_chk718 i_prm_oblgc_chk718(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[718])
);
prm_oblgc_chk719 i_prm_oblgc_chk719(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[719])
);
prm_oblgc_chk720 i_prm_oblgc_chk720(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[720])
);
prm_oblgc_chk721 i_prm_oblgc_chk721(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[721])
);
prm_oblgc_chk722 i_prm_oblgc_chk722(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[722])
);
prm_oblgc_chk723 i_prm_oblgc_chk723(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[723])
);
prm_oblgc_chk724 i_prm_oblgc_chk724(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[724])
);
prm_oblgc_chk725 i_prm_oblgc_chk725(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[725])
);
prm_oblgc_chk726 i_prm_oblgc_chk726(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[726])
);
prm_oblgc_chk727 i_prm_oblgc_chk727(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[727])
);
prm_oblgc_chk728 i_prm_oblgc_chk728(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[728])
);
prm_oblgc_chk729 i_prm_oblgc_chk729(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[729])
);
prm_oblgc_chk730 i_prm_oblgc_chk730(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[730])
);
prm_oblgc_chk731 i_prm_oblgc_chk731(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[731])
);
prm_oblgc_chk732 i_prm_oblgc_chk732(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[732])
);
prm_oblgc_chk733 i_prm_oblgc_chk733(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[733])
);
prm_oblgc_chk734 i_prm_oblgc_chk734(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[734])
);
prm_oblgc_chk735 i_prm_oblgc_chk735(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[735])
);
prm_oblgc_chk736 i_prm_oblgc_chk736(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[736])
);
prm_oblgc_chk737 i_prm_oblgc_chk737(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[737])
);
prm_oblgc_chk738 i_prm_oblgc_chk738(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[738])
);
prm_oblgc_chk739 i_prm_oblgc_chk739(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[739])
);
prm_oblgc_chk740 i_prm_oblgc_chk740(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[740])
);
prm_oblgc_chk741 i_prm_oblgc_chk741(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[741])
);
prm_oblgc_chk742 i_prm_oblgc_chk742(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[742])
);
prm_oblgc_chk743 i_prm_oblgc_chk743(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[743])
);
prm_oblgc_chk744 i_prm_oblgc_chk744(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[744])
);
prm_oblgc_chk745 i_prm_oblgc_chk745(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[745])
);
prm_oblgc_chk746 i_prm_oblgc_chk746(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[746])
);
prm_oblgc_chk747 i_prm_oblgc_chk747(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[747])
);
prm_oblgc_chk748 i_prm_oblgc_chk748(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[748])
);
prm_oblgc_chk749 i_prm_oblgc_chk749(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[749])
);
prm_oblgc_chk750 i_prm_oblgc_chk750(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[750])
);
prm_oblgc_chk751 i_prm_oblgc_chk751(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[751])
);
prm_oblgc_chk752 i_prm_oblgc_chk752(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[752])
);
prm_oblgc_chk753 i_prm_oblgc_chk753(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[753])
);
prm_oblgc_chk754 i_prm_oblgc_chk754(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[754])
);
prm_oblgc_chk755 i_prm_oblgc_chk755(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[755])
);
prm_oblgc_chk756 i_prm_oblgc_chk756(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[756])
);
prm_oblgc_chk757 i_prm_oblgc_chk757(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[757])
);
prm_oblgc_chk758 i_prm_oblgc_chk758(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[758])
);
prm_oblgc_chk759 i_prm_oblgc_chk759(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[759])
);
prm_oblgc_chk760 i_prm_oblgc_chk760(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[760])
);
prm_oblgc_chk761 i_prm_oblgc_chk761(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[761])
);
prm_oblgc_chk762 i_prm_oblgc_chk762(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[762])
);
prm_oblgc_chk763 i_prm_oblgc_chk763(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[763])
);
prm_oblgc_chk764 i_prm_oblgc_chk764(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[764])
);
prm_oblgc_chk765 i_prm_oblgc_chk765(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[765])
);
prm_oblgc_chk766 i_prm_oblgc_chk766(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[766])
);
prm_oblgc_chk767 i_prm_oblgc_chk767(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[767])
);
prm_oblgc_chk768 i_prm_oblgc_chk768(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[768])
);
prm_oblgc_chk769 i_prm_oblgc_chk769(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[769])
);
prm_oblgc_chk770 i_prm_oblgc_chk770(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[770])
);
prm_oblgc_chk771 i_prm_oblgc_chk771(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[771])
);
prm_oblgc_chk772 i_prm_oblgc_chk772(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[772])
);
prm_oblgc_chk773 i_prm_oblgc_chk773(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[773])
);
prm_oblgc_chk774 i_prm_oblgc_chk774(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[774])
);
prm_oblgc_chk775 i_prm_oblgc_chk775(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[775])
);
prm_oblgc_chk776 i_prm_oblgc_chk776(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[776])
);
prm_oblgc_chk777 i_prm_oblgc_chk777(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[777])
);
prm_oblgc_chk778 i_prm_oblgc_chk778(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[778])
);
prm_oblgc_chk779 i_prm_oblgc_chk779(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[779])
);
prm_oblgc_chk780 i_prm_oblgc_chk780(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[780])
);
prm_oblgc_chk781 i_prm_oblgc_chk781(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[781])
);
prm_oblgc_chk782 i_prm_oblgc_chk782(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[782])
);
prm_oblgc_chk783 i_prm_oblgc_chk783(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[783])
);
prm_oblgc_chk784 i_prm_oblgc_chk784(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[784])
);
prm_oblgc_chk785 i_prm_oblgc_chk785(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[785])
);
prm_oblgc_chk786 i_prm_oblgc_chk786(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[786])
);
prm_oblgc_chk787 i_prm_oblgc_chk787(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[787])
);
prm_oblgc_chk788 i_prm_oblgc_chk788(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[788])
);
prm_oblgc_chk789 i_prm_oblgc_chk789(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[789])
);
prm_oblgc_chk790 i_prm_oblgc_chk790(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[790])
);
prm_oblgc_chk791 i_prm_oblgc_chk791(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[791])
);
prm_oblgc_chk792 i_prm_oblgc_chk792(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[792])
);
prm_oblgc_chk793 i_prm_oblgc_chk793(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[793])
);
prm_oblgc_chk794 i_prm_oblgc_chk794(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[794])
);
prm_oblgc_chk795 i_prm_oblgc_chk795(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[795])
);
prm_oblgc_chk796 i_prm_oblgc_chk796(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[796])
);
prm_oblgc_chk797 i_prm_oblgc_chk797(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[797])
);
prm_oblgc_chk798 i_prm_oblgc_chk798(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[798])
);
prm_oblgc_chk799 i_prm_oblgc_chk799(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[799])
);
prm_oblgc_chk800 i_prm_oblgc_chk800(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[800])
);
prm_oblgc_chk801 i_prm_oblgc_chk801(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[801])
);
prm_oblgc_chk802 i_prm_oblgc_chk802(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[802])
);
prm_oblgc_chk803 i_prm_oblgc_chk803(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[803])
);
prm_oblgc_chk804 i_prm_oblgc_chk804(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[804])
);
prm_oblgc_chk805 i_prm_oblgc_chk805(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[805])
);
prm_oblgc_chk806 i_prm_oblgc_chk806(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[806])
);
prm_oblgc_chk807 i_prm_oblgc_chk807(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[807])
);
prm_oblgc_chk808 i_prm_oblgc_chk808(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[808])
);
prm_oblgc_chk809 i_prm_oblgc_chk809(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[809])
);
prm_oblgc_chk810 i_prm_oblgc_chk810(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[810])
);
prm_oblgc_chk811 i_prm_oblgc_chk811(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[811])
);
prm_oblgc_chk812 i_prm_oblgc_chk812(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[812])
);
prm_oblgc_chk813 i_prm_oblgc_chk813(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[813])
);
prm_oblgc_chk814 i_prm_oblgc_chk814(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[814])
);
prm_oblgc_chk815 i_prm_oblgc_chk815(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[815])
);
prm_oblgc_chk816 i_prm_oblgc_chk816(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[816])
);
prm_oblgc_chk817 i_prm_oblgc_chk817(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[817])
);
prm_oblgc_chk818 i_prm_oblgc_chk818(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[818])
);
prm_oblgc_chk819 i_prm_oblgc_chk819(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[819])
);
prm_oblgc_chk820 i_prm_oblgc_chk820(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[820])
);
prm_oblgc_chk821 i_prm_oblgc_chk821(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[821])
);
prm_oblgc_chk822 i_prm_oblgc_chk822(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[822])
);
prm_oblgc_chk823 i_prm_oblgc_chk823(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[823])
);
prm_oblgc_chk824 i_prm_oblgc_chk824(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[824])
);
prm_oblgc_chk825 i_prm_oblgc_chk825(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[825])
);
prm_oblgc_chk826 i_prm_oblgc_chk826(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[826])
);
prm_oblgc_chk827 i_prm_oblgc_chk827(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[827])
);
prm_oblgc_chk828 i_prm_oblgc_chk828(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[828])
);
prm_oblgc_chk829 i_prm_oblgc_chk829(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[829])
);
prm_oblgc_chk830 i_prm_oblgc_chk830(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[830])
);
prm_oblgc_chk831 i_prm_oblgc_chk831(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[831])
);
prm_oblgc_chk832 i_prm_oblgc_chk832(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[832])
);
prm_oblgc_chk833 i_prm_oblgc_chk833(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[833])
);
prm_oblgc_chk834 i_prm_oblgc_chk834(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[834])
);
prm_oblgc_chk835 i_prm_oblgc_chk835(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[835])
);
prm_oblgc_chk836 i_prm_oblgc_chk836(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[836])
);
prm_oblgc_chk837 i_prm_oblgc_chk837(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[837])
);
prm_oblgc_chk838 i_prm_oblgc_chk838(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[838])
);
prm_oblgc_chk839 i_prm_oblgc_chk839(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[839])
);
prm_oblgc_chk840 i_prm_oblgc_chk840(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[840])
);
prm_oblgc_chk841 i_prm_oblgc_chk841(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[841])
);
prm_oblgc_chk842 i_prm_oblgc_chk842(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[842])
);
prm_oblgc_chk843 i_prm_oblgc_chk843(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[843])
);
prm_oblgc_chk844 i_prm_oblgc_chk844(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[844])
);
prm_oblgc_chk845 i_prm_oblgc_chk845(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[845])
);
prm_oblgc_chk846 i_prm_oblgc_chk846(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[846])
);
prm_oblgc_chk847 i_prm_oblgc_chk847(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[847])
);
prm_oblgc_chk848 i_prm_oblgc_chk848(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[848])
);
prm_oblgc_chk849 i_prm_oblgc_chk849(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[849])
);
prm_oblgc_chk850 i_prm_oblgc_chk850(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[850])
);
prm_oblgc_chk851 i_prm_oblgc_chk851(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[851])
);
prm_oblgc_chk852 i_prm_oblgc_chk852(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[852])
);
prm_oblgc_chk853 i_prm_oblgc_chk853(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[853])
);
prm_oblgc_chk854 i_prm_oblgc_chk854(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[854])
);
prm_oblgc_chk855 i_prm_oblgc_chk855(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[855])
);
prm_oblgc_chk856 i_prm_oblgc_chk856(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[856])
);
prm_oblgc_chk857 i_prm_oblgc_chk857(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[857])
);
prm_oblgc_chk858 i_prm_oblgc_chk858(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[858])
);
prm_oblgc_chk859 i_prm_oblgc_chk859(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[859])
);
prm_oblgc_chk860 i_prm_oblgc_chk860(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[860])
);
prm_oblgc_chk861 i_prm_oblgc_chk861(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[861])
);
prm_oblgc_chk862 i_prm_oblgc_chk862(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[862])
);
prm_oblgc_chk863 i_prm_oblgc_chk863(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[863])
);
prm_oblgc_chk864 i_prm_oblgc_chk864(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[864])
);
prm_oblgc_chk865 i_prm_oblgc_chk865(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[865])
);
prm_oblgc_chk866 i_prm_oblgc_chk866(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[866])
);
prm_oblgc_chk867 i_prm_oblgc_chk867(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[867])
);
prm_oblgc_chk868 i_prm_oblgc_chk868(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[868])
);
prm_oblgc_chk869 i_prm_oblgc_chk869(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[869])
);
prm_oblgc_chk870 i_prm_oblgc_chk870(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[870])
);
prm_oblgc_chk871 i_prm_oblgc_chk871(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[871])
);
prm_oblgc_chk872 i_prm_oblgc_chk872(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[872])
);
prm_oblgc_chk873 i_prm_oblgc_chk873(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[873])
);
prm_oblgc_chk874 i_prm_oblgc_chk874(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[874])
);
prm_oblgc_chk875 i_prm_oblgc_chk875(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[875])
);
prm_oblgc_chk876 i_prm_oblgc_chk876(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[876])
);
prm_oblgc_chk877 i_prm_oblgc_chk877(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[877])
);
prm_oblgc_chk878 i_prm_oblgc_chk878(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[878])
);
prm_oblgc_chk879 i_prm_oblgc_chk879(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[879])
);
prm_oblgc_chk880 i_prm_oblgc_chk880(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[880])
);
prm_oblgc_chk881 i_prm_oblgc_chk881(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[881])
);
prm_oblgc_chk882 i_prm_oblgc_chk882(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[882])
);
prm_oblgc_chk883 i_prm_oblgc_chk883(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[883])
);
prm_oblgc_chk884 i_prm_oblgc_chk884(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[884])
);
prm_oblgc_chk885 i_prm_oblgc_chk885(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[885])
);
prm_oblgc_chk886 i_prm_oblgc_chk886(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[886])
);
prm_oblgc_chk887 i_prm_oblgc_chk887(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[887])
);
prm_oblgc_chk888 i_prm_oblgc_chk888(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[888])
);
prm_oblgc_chk889 i_prm_oblgc_chk889(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[889])
);
prm_oblgc_chk890 i_prm_oblgc_chk890(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[890])
);
prm_oblgc_chk891 i_prm_oblgc_chk891(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[891])
);
prm_oblgc_chk892 i_prm_oblgc_chk892(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[892])
);
prm_oblgc_chk893 i_prm_oblgc_chk893(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[893])
);
prm_oblgc_chk894 i_prm_oblgc_chk894(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[894])
);
prm_oblgc_chk895 i_prm_oblgc_chk895(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[895])
);
prm_oblgc_chk896 i_prm_oblgc_chk896(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[896])
);
prm_oblgc_chk897 i_prm_oblgc_chk897(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[897])
);
prm_oblgc_chk898 i_prm_oblgc_chk898(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[898])
);
prm_oblgc_chk899 i_prm_oblgc_chk899(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[899])
);
prm_oblgc_chk900 i_prm_oblgc_chk900(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[900])
);
prm_oblgc_chk901 i_prm_oblgc_chk901(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[901])
);
prm_oblgc_chk902 i_prm_oblgc_chk902(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[902])
);
prm_oblgc_chk903 i_prm_oblgc_chk903(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[903])
);
prm_oblgc_chk904 i_prm_oblgc_chk904(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[904])
);
prm_oblgc_chk905 i_prm_oblgc_chk905(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[905])
);
prm_oblgc_chk906 i_prm_oblgc_chk906(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[906])
);
prm_oblgc_chk907 i_prm_oblgc_chk907(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[907])
);
prm_oblgc_chk908 i_prm_oblgc_chk908(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[908])
);
prm_oblgc_chk909 i_prm_oblgc_chk909(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[909])
);
prm_oblgc_chk910 i_prm_oblgc_chk910(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[910])
);
prm_oblgc_chk911 i_prm_oblgc_chk911(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[911])
);
prm_oblgc_chk912 i_prm_oblgc_chk912(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[912])
);
prm_oblgc_chk913 i_prm_oblgc_chk913(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[913])
);
prm_oblgc_chk914 i_prm_oblgc_chk914(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[914])
);
prm_oblgc_chk915 i_prm_oblgc_chk915(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[915])
);
prm_oblgc_chk916 i_prm_oblgc_chk916(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[916])
);
prm_oblgc_chk917 i_prm_oblgc_chk917(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[917])
);
prm_oblgc_chk918 i_prm_oblgc_chk918(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[918])
);
prm_oblgc_chk919 i_prm_oblgc_chk919(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[919])
);
prm_oblgc_chk920 i_prm_oblgc_chk920(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[920])
);
prm_oblgc_chk921 i_prm_oblgc_chk921(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[921])
);
prm_oblgc_chk922 i_prm_oblgc_chk922(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[922])
);
prm_oblgc_chk923 i_prm_oblgc_chk923(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[923])
);
prm_oblgc_chk924 i_prm_oblgc_chk924(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[924])
);
prm_oblgc_chk925 i_prm_oblgc_chk925(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[925])
);
prm_oblgc_chk926 i_prm_oblgc_chk926(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[926])
);
prm_oblgc_chk927 i_prm_oblgc_chk927(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[927])
);
prm_oblgc_chk928 i_prm_oblgc_chk928(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[928])
);
prm_oblgc_chk929 i_prm_oblgc_chk929(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[929])
);
prm_oblgc_chk930 i_prm_oblgc_chk930(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[930])
);
prm_oblgc_chk931 i_prm_oblgc_chk931(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[931])
);
prm_oblgc_chk932 i_prm_oblgc_chk932(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[932])
);
prm_oblgc_chk933 i_prm_oblgc_chk933(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[933])
);
prm_oblgc_chk934 i_prm_oblgc_chk934(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[934])
);
prm_oblgc_chk935 i_prm_oblgc_chk935(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[935])
);
prm_oblgc_chk936 i_prm_oblgc_chk936(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[936])
);
prm_oblgc_chk937 i_prm_oblgc_chk937(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[937])
);
prm_oblgc_chk938 i_prm_oblgc_chk938(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[938])
);
prm_oblgc_chk939 i_prm_oblgc_chk939(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[939])
);
prm_oblgc_chk940 i_prm_oblgc_chk940(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[940])
);
prm_oblgc_chk941 i_prm_oblgc_chk941(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[941])
);
prm_oblgc_chk942 i_prm_oblgc_chk942(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[942])
);
prm_oblgc_chk943 i_prm_oblgc_chk943(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[943])
);
prm_oblgc_chk944 i_prm_oblgc_chk944(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[944])
);
prm_oblgc_chk945 i_prm_oblgc_chk945(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[945])
);
prm_oblgc_chk946 i_prm_oblgc_chk946(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[946])
);
prm_oblgc_chk947 i_prm_oblgc_chk947(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[947])
);
prm_oblgc_chk948 i_prm_oblgc_chk948(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[948])
);
prm_oblgc_chk949 i_prm_oblgc_chk949(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[949])
);
prm_oblgc_chk950 i_prm_oblgc_chk950(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[950])
);
prm_oblgc_chk951 i_prm_oblgc_chk951(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[951])
);
prm_oblgc_chk952 i_prm_oblgc_chk952(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[952])
);
prm_oblgc_chk953 i_prm_oblgc_chk953(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[953])
);
prm_oblgc_chk954 i_prm_oblgc_chk954(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[954])
);
prm_oblgc_chk955 i_prm_oblgc_chk955(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[955])
);
prm_oblgc_chk956 i_prm_oblgc_chk956(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[956])
);
prm_oblgc_chk957 i_prm_oblgc_chk957(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[957])
);
prm_oblgc_chk958 i_prm_oblgc_chk958(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[958])
);
prm_oblgc_chk959 i_prm_oblgc_chk959(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[959])
);
prm_oblgc_chk960 i_prm_oblgc_chk960(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[960])
);
prm_oblgc_chk961 i_prm_oblgc_chk961(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[961])
);
prm_oblgc_chk962 i_prm_oblgc_chk962(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[962])
);
prm_oblgc_chk963 i_prm_oblgc_chk963(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[963])
);
prm_oblgc_chk964 i_prm_oblgc_chk964(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[964])
);
prm_oblgc_chk965 i_prm_oblgc_chk965(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[965])
);
prm_oblgc_chk966 i_prm_oblgc_chk966(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[966])
);
prm_oblgc_chk967 i_prm_oblgc_chk967(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[967])
);
prm_oblgc_chk968 i_prm_oblgc_chk968(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[968])
);
prm_oblgc_chk969 i_prm_oblgc_chk969(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[969])
);
prm_oblgc_chk970 i_prm_oblgc_chk970(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[970])
);
prm_oblgc_chk971 i_prm_oblgc_chk971(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[971])
);
prm_oblgc_chk972 i_prm_oblgc_chk972(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[972])
);
prm_oblgc_chk973 i_prm_oblgc_chk973(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[973])
);
prm_oblgc_chk974 i_prm_oblgc_chk974(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[974])
);
prm_oblgc_chk975 i_prm_oblgc_chk975(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[975])
);
prm_oblgc_chk976 i_prm_oblgc_chk976(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[976])
);
prm_oblgc_chk977 i_prm_oblgc_chk977(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[977])
);
prm_oblgc_chk978 i_prm_oblgc_chk978(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[978])
);
prm_oblgc_chk979 i_prm_oblgc_chk979(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[979])
);
prm_oblgc_chk980 i_prm_oblgc_chk980(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[980])
);
prm_oblgc_chk981 i_prm_oblgc_chk981(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[981])
);
prm_oblgc_chk982 i_prm_oblgc_chk982(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[982])
);
prm_oblgc_chk983 i_prm_oblgc_chk983(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[983])
);
prm_oblgc_chk984 i_prm_oblgc_chk984(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[984])
);
prm_oblgc_chk985 i_prm_oblgc_chk985(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[985])
);
prm_oblgc_chk986 i_prm_oblgc_chk986(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[986])
);
prm_oblgc_chk987 i_prm_oblgc_chk987(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[987])
);
prm_oblgc_chk988 i_prm_oblgc_chk988(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[988])
);
prm_oblgc_chk989 i_prm_oblgc_chk989(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[989])
);
prm_oblgc_chk990 i_prm_oblgc_chk990(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[990])
);
prm_oblgc_chk991 i_prm_oblgc_chk991(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[991])
);
prm_oblgc_chk992 i_prm_oblgc_chk992(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[992])
);
prm_oblgc_chk993 i_prm_oblgc_chk993(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[993])
);
prm_oblgc_chk994 i_prm_oblgc_chk994(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[994])
);
prm_oblgc_chk995 i_prm_oblgc_chk995(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[995])
);
prm_oblgc_chk996 i_prm_oblgc_chk996(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[996])
);
prm_oblgc_chk997 i_prm_oblgc_chk997(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[997])
);
prm_oblgc_chk998 i_prm_oblgc_chk998(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[998])
);
prm_oblgc_chk999 i_prm_oblgc_chk999(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[999])
);
prm_oblgc_chk1000 i_prm_oblgc_chk1000(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1000])
);
prm_oblgc_chk1001 i_prm_oblgc_chk1001(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1001])
);
prm_oblgc_chk1002 i_prm_oblgc_chk1002(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1002])
);
prm_oblgc_chk1003 i_prm_oblgc_chk1003(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1003])
);
prm_oblgc_chk1004 i_prm_oblgc_chk1004(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1004])
);
prm_oblgc_chk1005 i_prm_oblgc_chk1005(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1005])
);
prm_oblgc_chk1006 i_prm_oblgc_chk1006(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1006])
);
prm_oblgc_chk1007 i_prm_oblgc_chk1007(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1007])
);
prm_oblgc_chk1008 i_prm_oblgc_chk1008(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1008])
);
prm_oblgc_chk1009 i_prm_oblgc_chk1009(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1009])
);
prm_oblgc_chk1010 i_prm_oblgc_chk1010(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1010])
);
prm_oblgc_chk1011 i_prm_oblgc_chk1011(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1011])
);
prm_oblgc_chk1012 i_prm_oblgc_chk1012(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1012])
);
prm_oblgc_chk1013 i_prm_oblgc_chk1013(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1013])
);
prm_oblgc_chk1014 i_prm_oblgc_chk1014(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1014])
);
prm_oblgc_chk1015 i_prm_oblgc_chk1015(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1015])
);
prm_oblgc_chk1016 i_prm_oblgc_chk1016(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1016])
);
prm_oblgc_chk1017 i_prm_oblgc_chk1017(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1017])
);
prm_oblgc_chk1018 i_prm_oblgc_chk1018(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1018])
);
prm_oblgc_chk1019 i_prm_oblgc_chk1019(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1019])
);
prm_oblgc_chk1020 i_prm_oblgc_chk1020(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1020])
);
prm_oblgc_chk1021 i_prm_oblgc_chk1021(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1021])
);
prm_oblgc_chk1022 i_prm_oblgc_chk1022(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1022])
);
prm_oblgc_chk1023 i_prm_oblgc_chk1023(
.A(A),
.B(B),
.C(C),
.D(D),
.E(E),
.F(F),
.G(G),
.H(H),
.I(I),
.J(J),
.K(K),
.L(L),
.M(M),
.N(N),
.O(O),
.edge_mask(edge_mask[1023])
);
endmodule
